`timescale 1ns / 1ps  

module testbench ();
	
	reg[15:0] in1, in2;
	reg sel;
	wire[15:0] out;

	mux21 u (in1, in2, sel, out);

initial
begin
	in1 = 0;
	in2 = 0;
	sel = 0;
	#50 in1 = 1;
	in2 = 2;
	sel = 0;
	#50 sel = 1;
	#50;
end

endmodule
