`timescale 1ns / 1ps

module testbench ();
  parameter ADDR_BIT = 6;
  parameter DATA_BIT = 16;
  parameter N = 256;
  parameter n = 8;
  parameter MEM_HEIGHT = N / 4;

  
  /* all the input data is stored here */  
  //reg [DATA_BIT * MEM_HEIGHT * 4 - 1 : 0] input_data;
  parameter [DATA_BIT - 1 : 0] input_data[0 : N - 1] = '{16'b0, {15'b0, 1'b1}, {14'b0, 2'b10}, {14'b0, 2'b11}, {13'b0, 3'b100}, {13'b0, 3'b101}, {13'b0, 3'b110}, {13'b0, 3'b111}, {12'b0, 4'b1000}, {12'b0, 4'b1001}, {12'b0, 4'b1010}, {12'b0, 4'b1011}, {12'b0, 4'b1100}, {12'b0, 4'b1101}, {12'b0, 4'b1110}, {12'b0, 4'b1111}, {11'b0, 5'b10000}, {11'b0, 5'b10001}, {11'b0, 5'b10010}, {11'b0, 5'b10011}, {11'b0, 5'b10100}, {11'b0, 5'b10101}, {11'b0, 5'b10110}, {11'b0, 5'b10111}, {11'b0, 5'b11000}, {11'b0, 5'b11001}, {11'b0, 5'b11010}, {11'b0, 5'b11011}, {11'b0, 5'b11100}, {11'b0, 5'b11101}, {11'b0, 5'b11110}, {11'b0,5'b11111}, 16'b0, {15'b0, 1'b1}, {14'b0, 2'b10}, {14'b0, 2'b11}, {13'b0, 3'b100}, {13'b0, 3'b101}, {13'b0, 3'b110}, {13'b0, 3'b111}, {12'b0, 4'b1000}, {12'b0, 4'b1001}, {12'b0, 4'b1010}, {12'b0, 4'b1011}, {12'b0, 4'b1100}, {12'b0, 4'b1101}, {12'b0, 4'b1110}, {12'b0, 4'b1111}, {11'b0, 5'b10000}, {11'b0, 5'b10001}, {11'b0, 5'b10010}, {11'b0, 5'b10011}, {11'b0, 5'b10100}, {11'b0, 5'b10101}, {11'b0, 5'b10110}, {11'b0, 5'b10111}, {11'b0, 5'b11000}, {11'b0, 5'b11001}, {11'b0, 5'b11010}, {11'b0, 5'b11011}, {11'b0, 5'b11100}, {11'b0, 5'b11101}, {11'b0, 5'b11110}, {11'b0,5'b11111},16'b0, {15'b0, 1'b1}, {14'b0, 2'b10}, {14'b0, 2'b11}, {13'b0, 3'b100}, {13'b0, 3'b101}, {13'b0, 3'b110}, {13'b0, 3'b111}, {12'b0, 4'b1000}, {12'b0, 4'b1001}, {12'b0, 4'b1010}, {12'b0, 4'b1011}, {12'b0, 4'b1100}, {12'b0, 4'b1101}, {12'b0, 4'b1110}, {12'b0, 4'b1111}, {11'b0, 5'b10000}, {11'b0, 5'b10001}, {11'b0, 5'b10010}, {11'b0, 5'b10011}, {11'b0, 5'b10100}, {11'b0, 5'b10101}, {11'b0, 5'b10110}, {11'b0, 5'b10111}, {11'b0, 5'b11000}, {11'b0, 5'b11001}, {11'b0, 5'b11010}, {11'b0, 5'b11011}, {11'b0, 5'b11100}, {11'b0, 5'b11101}, {11'b0, 5'b11110}, {11'b0,5'b11111},16'b0, {15'b0, 1'b1}, {14'b0, 2'b10}, {14'b0, 2'b11}, {13'b0, 3'b100}, {13'b0, 3'b101}, {13'b0, 3'b110}, {13'b0, 3'b111}, {12'b0, 4'b1000}, {12'b0, 4'b1001}, {12'b0, 4'b1010}, {12'b0, 4'b1011}, {12'b0, 4'b1100}, {12'b0, 4'b1101}, {12'b0, 4'b1110}, {12'b0, 4'b1111}, {11'b0, 5'b10000}, {11'b0, 5'b10001}, {11'b0, 5'b10010}, {11'b0, 5'b10011}, {11'b0, 5'b10100}, {11'b0, 5'b10101}, {11'b0, 5'b10110}, {11'b0, 5'b10111}, {11'b0, 5'b11000}, {11'b0, 5'b11001}, {11'b0, 5'b11010}, {11'b0, 5'b11011}, {11'b0, 5'b11100}, {11'b0, 5'b11101}, {11'b0, 5'b11110}, {11'b0,5'b11111}, 16'b0, {15'b0, 1'b1}, {14'b0, 2'b10}, {14'b0, 2'b11}, {13'b0, 3'b100}, {13'b0, 3'b101}, {13'b0, 3'b110}, {13'b0, 3'b111}, {12'b0, 4'b1000}, {12'b0, 4'b1001}, {12'b0, 4'b1010}, {12'b0, 4'b1011}, {12'b0, 4'b1100}, {12'b0, 4'b1101}, {12'b0, 4'b1110}, {12'b0, 4'b1111}, {11'b0, 5'b10000}, {11'b0, 5'b10001}, {11'b0, 5'b10010}, {11'b0, 5'b10011}, {11'b0, 5'b10100}, {11'b0, 5'b10101}, {11'b0, 5'b10110}, {11'b0, 5'b10111}, {11'b0, 5'b11000}, {11'b0, 5'b11001}, {11'b0, 5'b11010}, {11'b0, 5'b11011}, {11'b0, 5'b11100}, {11'b0, 5'b11101}, {11'b0, 5'b11110}, {11'b0,5'b11111}, 16'b0, {15'b0, 1'b1}, {14'b0, 2'b10}, {14'b0, 2'b11}, {13'b0, 3'b100}, {13'b0, 3'b101}, {13'b0, 3'b110}, {13'b0, 3'b111}, {12'b0, 4'b1000}, {12'b0, 4'b1001}, {12'b0, 4'b1010}, {12'b0, 4'b1011}, {12'b0, 4'b1100}, {12'b0, 4'b1101}, {12'b0, 4'b1110}, {12'b0, 4'b1111}, {11'b0, 5'b10000}, {11'b0, 5'b10001}, {11'b0, 5'b10010}, {11'b0, 5'b10011}, {11'b0, 5'b10100}, {11'b0, 5'b10101}, {11'b0, 5'b10110}, {11'b0, 5'b10111}, {11'b0, 5'b11000}, {11'b0, 5'b11001}, {11'b0, 5'b11010}, {11'b0, 5'b11011}, {11'b0, 5'b11100}, {11'b0, 5'b11101}, {11'b0, 5'b11110}, {11'b0,5'b11111},16'b0, {15'b0, 1'b1}, {14'b0, 2'b10}, {14'b0, 2'b11}, {13'b0, 3'b100}, {13'b0, 3'b101}, {13'b0, 3'b110}, {13'b0, 3'b111}, {12'b0, 4'b1000}, {12'b0, 4'b1001}, {12'b0, 4'b1010}, {12'b0, 4'b1011}, {12'b0, 4'b1100}, {12'b0, 4'b1101}, {12'b0, 4'b1110}, {12'b0, 4'b1111}, {11'b0, 5'b10000}, {11'b0, 5'b10001}, {11'b0, 5'b10010}, {11'b0, 5'b10011}, {11'b0, 5'b10100}, {11'b0, 5'b10101}, {11'b0, 5'b10110}, {11'b0, 5'b10111}, {11'b0, 5'b11000}, {11'b0, 5'b11001}, {11'b0, 5'b11010}, {11'b0, 5'b11011}, {11'b0, 5'b11100}, {11'b0, 5'b11101}, {11'b0, 5'b11110}, {11'b0,5'b11111},16'b0, {15'b0, 1'b1}, {14'b0, 2'b10}, {14'b0, 2'b11}, {13'b0, 3'b100}, {13'b0, 3'b101}, {13'b0, 3'b110}, {13'b0, 3'b111}, {12'b0, 4'b1000}, {12'b0, 4'b1001}, {12'b0, 4'b1010}, {12'b0, 4'b1011}, {12'b0, 4'b1100}, {12'b0, 4'b1101}, {12'b0, 4'b1110}, {12'b0, 4'b1111}, {11'b0, 5'b10000}, {11'b0, 5'b10001}, {11'b0, 5'b10010}, {11'b0, 5'b10011}, {11'b0, 5'b10100}, {11'b0, 5'b10101}, {11'b0, 5'b10110}, {11'b0, 5'b10111}, {11'b0, 5'b11000}, {11'b0, 5'b11001}, {11'b0, 5'b11010}, {11'b0, 5'b11011}, {11'b0, 5'b11100}, {11'b0, 5'b11101}, {11'b0, 5'b11110}, {11'b0,5'b11111}};

  reg [DATA_BIT - 1 : 0] in0, in1, in2, in3, w_r, w_i;
  reg clk;
  reg rst;
  reg rst_top;
  wire [DATA_BIT - 1 : 0] mem0_i, mem1_i, mem2_i, mem3_i;
  wire [DATA_BIT - 1 : 0] mem0_o, mem1_o, mem2_o, mem3_o;
  wire [DATA_BIT - 1 : 0] mem0, mem1, mem2, mem3;
  reg [1 : 0] m12, m13;
  reg [ADDR_BIT * 4 - 1 : 0] addr_read, addr_write;
  reg [ADDR_BIT - 1 : 0] upcounter;
  reg bypass_en;
  //reg [ADDR_BIT - 1 : 0] read_s_index;
  //reg start;
  //reg rst;
  reg prepare_data;
  reg [DATA_BIT - 1 : 0] input_d0;
  reg [DATA_BIT - 1 : 0] input_d1;
  reg [DATA_BIT - 1 : 0] input_d2;
  reg [DATA_BIT - 1 : 0] input_d3;
  reg [3 : 0] stage;
  
  
  top_level tl(prepare_data, clk, rst_top, input_d0, input_d1, input_d2, input_d3, mem0_o, mem1_o, mem2_o, mem3_o);
 
  /* stage counter */
  always @(upcounter /*or prepare_data*/)
        if (upcounter == 6'b000000)
                stage = stage + 1;

  /* cycle counter for each stage */
  always @(posedge clk)
	if (rst)
		upcounter <= 0;
	else
		upcounter <= upcounter + 1;
	
  /* twiddle setup */


  /* load data control */
  always @(upcounter)
	begin
	if (prepare_data)
		begin
		input_d0 = input_data[upcounter];
                input_d1 = input_data[MEM_HEIGHT + upcounter];
                input_d2 = input_data[MEM_HEIGHT * 2 + upcounter];
                input_d3 = input_data[MEM_HEIGHT * 3 + upcounter];
		end
	end


  /* data input */
  

  initial begin
	clk = 1;
	rst = 1;
	rst_top = 1;
	#20
	rst = 0;
	rst_top = 1;
	upcounter = 6'b111111;
	prepare_data = 1;
	stage = 0;
	#640
	prepare_data = 0;
	rst_top = 0;	
			
	
    
  end

  always
    #5 clk = ~clk;

endmodule // testbench
